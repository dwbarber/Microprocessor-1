
class sequence_item extends uvm_sequence_item;
    //signals

    rand logic [3:0] a, b; //randomizeable inputs
    logic [4:0] sum; //output

endclass